module TEST_MUX (

	input [7:0] in,
	input sel,
	output [7:0] data_a,
	output [7:0] data_b
);

reg [7:0] o;

always@(*)
	begin
		case(sel)
		1'b0: o =
		
	end
endmodule
	
