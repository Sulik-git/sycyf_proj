module ADD_RSP_CHECK(
	
	input clk,
	input add_rsp,
	output next


);

reg next_local;

always@(posedge clk)begin

		next_local = 


end